module inverter (a,YINV);
input a;
output YINV;
assign YINV =~a;
endmodule